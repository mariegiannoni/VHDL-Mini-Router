library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.numeric_std.all;

---------
-- LUT --
---------

entity LUT is
	Port(
		lut_in : in std_logic_vector(6 downto 0);
		lut_out : out std_logic_vector(2 downto 0)
	);
end LUT;

architecture rtl of LUT is
signal lut_in_integer : integer range 0 to 127;
type lut_t is array (natural range<>) of std_logic_vector(2 downto 0);
constant lut : lut_t (0 to 127) := (
					"000",
					"001",
					"000",
					"001",
					"000",
					"001",
					"000",
					"001",
					"000",
					"001",
					"000",
					"001",
					"000",
					"001",
					"000",
					"001",
					"000",
					"001",
					"000",
					"001",
					"000",
					"001",
					"000",
					"001",
					"000",
					"001",
					"000",
					"001",
					"000",
					"001",
					"000",
					"001",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"101",
					"110",
					"110",
					"111",
					"100",
					"101",
					"101",
					"110",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"110",
					"111",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"100",
					"101",
					"101",
					"110",
					"110",
					"111",
					"100",
					"101",
					"101",
					"110"
				    );

begin
	-- we convert the 7 bits input in an integer from 0 to 127. 0 to  127 is the range of the 3 bits value in the look-up table.
	lut_in_integer <= TO_INTEGER(unsigned(lut_in));
	-- we retrive in the look-up table the element with the range previously computed
	lut_out <= lut(lut_in_integer);
end rtl;